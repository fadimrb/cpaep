module adder_tree #(
  /*automatically generates an adder tree, possibly pipelined, to add more than two numbers together*/

  parameter int ADDEND_WIDTH = 32,               // width of the addends
  parameter int OUT_SCALE = 0,                   // by how many bits to downscale the output
  parameter int OUT_WIDTH = 32,                  // the width of the output
  parameter int NB_ADDENDS = 4,                  // the number of addends to be summed
  parameter int NB_LEVELS_IN_PIPELINE_STAGE = 2  // after every this amount of levels of the adder tree, pipeline registers are added
  )
  (
  input logic clk, arst_n_in, // both of these can be left open if NB_LEVELS_IN_PIPELINE_STAGE > ceil(log2(NB_ADDENDS)), as then there is no pipelining
  input logic signed [ADDEND_WIDTH-1:0] addends[0:NB_ADDENDS-1],
  output logic signed [OUT_WIDTH-1:0] out
  );

  // every level of an adder tree divides the number of addends still to add by 2, so we need this many levels
  localparam NB_LEVELS = $clog2(NB_ADDENDS);
  localparam PSUM_WIDTH = OUT_WIDTH + OUT_SCALE; // higher significant bits will be thrown away at the end anyways

  // the partial sums (including inputs and unscaled output), passed between levels
  logic signed [PSUM_WIDTH-1:0] psums[0:NB_LEVELS][0:NB_ADDENDS-1]; // this is a rectangular matrix of psums, although only a triangle is needed.
                                                             // A triangle is much more complex though. So we just instantiate all these wires.
                                                             // Any synthesis tools would easily remove the redundant wires.

  assign psums[0] = addends;

  generate
    genvar level, a_in_level;
    //level 0 is just the inputs
    //so we start at level 1
    for (level = 1; level <= NB_LEVELS; level = level + 1) begin:level_loop
      //in every level, we loop over a counter that runs up to NB_ADDENDS so that we can set all the elements of psums
      //A part of these will be sums of psums of the previous level, generated by adders
      //then there is possibly a copy of a psum of the previous level, if there is an odd amount
      //the rest is filled with x's as they are useless signals.
      for (a_in_level = 0; a_in_level < NB_ADDENDS; a_in_level = a_in_level + 1) begin: a_in_level_loop
        logic signed [PSUM_WIDTH-1:0] unlatched_psum;
        if ((a_in_level) < ((NB_ADDENDS + ((1<<(level-1)) -1 )) / (1<<(level-1)))/2) begin: a_in_usefull_range
          // for these we need an adder
          adder #(.A_WIDTH(PSUM_WIDTH),
                  .B_WIDTH(PSUM_WIDTH),
                  .OUT_WIDTH(PSUM_WIDTH),
                  .OUT_SCALE(0))
                  adder_i
                  (.a(psums[level-1][a_in_level*2]),
                   .b(psums[level-1][a_in_level*2 +1]),
                   .out(unlatched_psum));
          // add pipeline registers if necessary at this stage
          if (level % NB_LEVELS_IN_PIPELINE_STAGE == 0) begin:if_with_pipeline
            register #(.WIDTH(PSUM_WIDTH), .RESET_VAL(0))
              pipeline_register_i
                (.clk(clk),
                 .arst_n_in(arst_n_in),
                 .din(unlatched_psum),
                 .qout(psums[level][a_in_level]),
                 .we(1'b1));
          end else begin:else_just_assign // else just assign unlatched output directly
            assign psums[level][a_in_level] = unlatched_psum;
          end


        end else if ((a_in_level+1)*2 == ((NB_ADDENDS + ((1<<(level-1)) -1 )) / (1<<(level-1)))+1) begin: odd_addend
          //We don't need an extra adder, but there is an odd addend left, we just pass this on to the next level
          assign unlatched_psum = psums[level-1][a_in_level*2];
          // add pipeline registers if necessary at this stage
          if (level % NB_LEVELS_IN_PIPELINE_STAGE == 0) begin:if_with_pipeline
            register #(.WIDTH(PSUM_WIDTH), .RESET_VAL(0))
              pipeline_register_i
                (.clk(clk),
                 .arst_n_in(arst_n_in),
                 .din(unlatched_psum),
                 .qout(psums[level][a_in_level]),
                 .we(1'b1));
          end else begin:else_just_assign // else just assign unlatched output directly
            assign psums[level][a_in_level] = unlatched_psum;
          end

        end else begin:a_outside_usefull_range
          //These signals are not necessary in this level (fall outside the triangle)
          assign psums[level][a_in_level] = 'x;
        end
      end
    end
  endgenerate

  //Finally, let's not forget the output scaling. 
  assign out = psums[NB_LEVELS][0] >>> OUT_SCALE;

endmodule
